magic
tech sky130A
magscale 1 2
timestamp 1729233261
<< nwell >>
rect -184 -877 814 1995
<< nsubdiff >>
rect -148 1925 -83 1959
rect 709 1925 778 1959
rect -148 1897 -114 1925
rect 744 1897 778 1925
rect -148 -807 -114 -745
rect 744 -807 778 -745
rect -148 -841 -83 -807
rect 709 -841 778 -807
<< nsubdiffcont >>
rect -83 1925 709 1959
rect -148 -745 -114 1897
rect 744 -745 778 1897
rect -83 -841 709 -807
<< poly >>
rect -64 1887 28 1903
rect -64 1853 -48 1887
rect -14 1853 28 1887
rect -64 1838 28 1853
rect -2 1818 28 1838
rect 602 1887 694 1903
rect 602 1853 644 1887
rect 678 1853 694 1887
rect 602 1838 694 1853
rect 602 1818 632 1838
rect -64 1193 28 1209
rect 86 1208 286 1310
rect -64 1159 -48 1193
rect -14 1159 28 1193
rect -64 1144 28 1159
rect -2 1124 28 1144
rect 602 1193 694 1209
rect 602 1159 644 1193
rect 678 1159 694 1193
rect 602 1144 694 1159
rect 602 1126 632 1144
rect -64 499 28 515
rect 86 514 544 616
rect -64 465 -48 499
rect -14 465 28 499
rect -64 450 28 465
rect -2 430 28 450
rect 602 499 694 515
rect 602 465 644 499
rect 678 465 694 499
rect 602 450 694 465
rect 602 430 632 450
rect 344 -180 544 -78
rect 602 -183 694 -167
rect 602 -217 644 -183
rect 678 -217 694 -183
rect 602 -232 694 -217
rect 602 -250 632 -232
rect -2 -720 28 -702
rect -64 -735 28 -720
rect -64 -769 -48 -735
rect -14 -769 28 -735
rect -64 -785 28 -769
<< polycont >>
rect -48 1853 -14 1887
rect 644 1853 678 1887
rect -48 1159 -14 1193
rect 644 1159 678 1193
rect -48 465 -14 499
rect 644 465 678 499
rect 644 -217 678 -183
rect -48 -769 -14 -735
<< locali >>
rect -148 1925 -83 1959
rect 709 1925 778 1959
rect -148 1897 -114 1925
rect 744 1897 778 1925
rect -64 1853 -48 1887
rect -14 1853 2 1887
rect 628 1853 644 1887
rect 678 1853 694 1887
rect -48 1790 -14 1853
rect 644 1788 678 1853
rect -64 1159 -48 1193
rect -14 1159 2 1193
rect 628 1159 644 1193
rect 678 1159 694 1193
rect -48 1096 -14 1159
rect 644 1094 678 1159
rect -64 465 -48 499
rect -14 465 2 499
rect 628 465 644 499
rect 678 465 694 499
rect -48 402 -14 465
rect 644 402 678 465
rect 628 -217 644 -183
rect 678 -217 694 -183
rect -48 -290 -14 -275
rect 644 -291 678 -217
rect -48 -735 -14 -661
rect -148 -807 -114 -745
rect -64 -769 -48 -735
rect -14 -769 2 -735
rect 744 -807 778 -745
rect -148 -841 -83 -807
rect 709 -841 778 -807
<< viali >>
rect 644 1925 678 1959
rect -48 1853 -14 1887
rect 644 1853 678 1887
rect -48 1159 -14 1193
rect 644 1159 678 1193
rect -48 465 -14 499
rect 644 465 678 499
rect 644 -217 678 -183
rect -48 -769 -14 -735
rect -48 -841 -14 -807
<< metal1 >>
rect 632 1959 690 1965
rect 632 1925 644 1959
rect 678 1925 690 1959
rect -60 1887 -2 1893
rect -60 1853 -48 1887
rect -14 1853 -2 1887
rect -60 1847 -2 1853
rect 632 1887 690 1925
rect 632 1853 644 1887
rect 678 1853 690 1887
rect 632 1847 690 1853
rect -54 1806 -8 1847
rect 638 1806 684 1847
rect -54 1794 80 1806
rect -66 1418 -56 1794
rect -4 1418 80 1794
rect -54 1406 80 1418
rect 298 1364 332 1418
rect 550 1406 684 1806
rect 550 1364 596 1406
rect 298 1320 596 1364
rect -60 1193 -2 1199
rect -60 1159 -48 1193
rect -14 1159 -2 1193
rect -60 1153 -2 1159
rect -54 1112 -8 1153
rect -54 1100 80 1112
rect -54 724 32 1100
rect 84 724 94 1100
rect -54 712 80 724
rect -60 499 -2 505
rect -60 465 -48 499
rect -14 465 -2 499
rect 54 481 134 502
rect -60 459 -2 465
rect 38 462 134 481
rect -54 418 -8 459
rect 38 418 76 462
rect -54 18 80 418
rect 298 -190 332 1320
rect 632 1193 690 1199
rect 632 1159 644 1193
rect 678 1159 690 1193
rect 632 1153 690 1159
rect 636 1112 688 1153
rect 550 1084 688 1112
rect 550 712 684 1084
rect 554 668 594 712
rect 498 628 594 668
rect 632 499 690 505
rect 632 465 644 499
rect 678 465 690 499
rect 632 459 690 465
rect 638 418 684 459
rect 550 406 684 418
rect 538 30 548 406
rect 600 30 684 406
rect 550 18 684 30
rect 34 -234 332 -190
rect 632 -183 690 -167
rect 632 -217 644 -183
rect 678 -217 690 -183
rect 632 -223 690 -217
rect -54 -276 -8 -275
rect 34 -276 80 -234
rect -54 -676 80 -276
rect 298 -288 332 -234
rect 636 -276 688 -223
rect 550 -288 688 -276
rect 550 -664 636 -288
rect 688 -664 698 -288
rect 550 -676 684 -664
rect -54 -729 -8 -676
rect -60 -735 -2 -729
rect -60 -769 -48 -735
rect -14 -769 -2 -735
rect -60 -807 -2 -769
rect -60 -841 -48 -807
rect -14 -841 -2 -807
rect -60 -847 -2 -841
<< via1 >>
rect -56 1418 -4 1794
rect 32 724 84 1100
rect 548 30 600 406
rect 636 -664 688 -288
<< metal2 >>
rect -56 1794 -4 1804
rect -56 1312 -4 1418
rect -58 1302 -2 1312
rect -58 1224 -2 1234
rect 628 1296 692 1306
rect 628 1230 692 1240
rect -56 -90 -4 1224
rect 32 1100 84 1110
rect 32 596 84 724
rect 32 542 600 596
rect 548 406 600 542
rect 548 20 600 30
rect 636 -90 688 1230
rect -58 -100 -2 -90
rect -58 -166 -2 -156
rect 634 -100 690 -90
rect 634 -166 690 -156
rect 636 -288 688 -166
rect 636 -674 688 -664
<< via2 >>
rect -58 1234 -2 1302
rect 628 1240 692 1296
rect -58 -156 -2 -100
rect 634 -156 690 -100
<< metal3 >>
rect -68 1302 8 1307
rect -68 1234 -58 1302
rect -2 1296 702 1302
rect -2 1240 628 1296
rect 692 1240 702 1296
rect -2 1234 702 1240
rect -68 1229 8 1234
rect -68 -100 700 -94
rect -68 -156 -58 -100
rect -2 -156 634 -100
rect 690 -156 700 -100
rect -68 -162 700 -156
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_0
timestamp 1729233261
transform 1 0 13 0 1 218
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_1
timestamp 1729233261
transform 1 0 13 0 1 -476
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_2
timestamp 1729233261
transform 1 0 617 0 1 -476
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_3
timestamp 1729233261
transform 1 0 617 0 1 218
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_4
timestamp 1729233261
transform 1 0 617 0 1 912
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_5
timestamp 1729233261
transform 1 0 617 0 1 1606
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_6
timestamp 1729233261
transform 1 0 13 0 1 1606
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_7
timestamp 1729233261
transform 1 0 13 0 1 912
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_0
timestamp 1729233261
transform 1 0 315 0 1 1606
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_1
timestamp 1729233261
transform 1 0 315 0 1 912
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_2
timestamp 1729233261
transform 1 0 315 0 1 218
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_3
timestamp 1729233261
transform 1 0 315 0 1 -476
box -323 -300 323 300
<< labels >>
flabel metal1 658 1917 658 1917 0 FreeSans 160 0 0 0 VDD
port 0 nsew
flabel metal2 662 606 662 606 0 FreeSans 160 0 0 0 D5
port 1 nsew
flabel metal1 572 659 572 659 0 FreeSans 160 0 0 0 D2
port 2 nsew
flabel metal2 59 625 59 625 0 FreeSans 160 0 0 0 D1
port 3 nsew
<< end >>
