magic
tech sky130A
magscale 1 2
timestamp 1729213131
<< nwell >>
rect -306 -578 1411 494
<< nsubdiff >>
rect -270 424 -201 458
rect 1309 424 1375 458
rect -270 389 -236 424
rect -270 -508 -236 -483
rect 1341 389 1375 424
rect 1341 -508 1375 -483
rect -270 -542 -201 -508
rect 1309 -542 1375 -508
<< nsubdiffcont >>
rect -201 424 1309 458
rect -270 -483 -236 389
rect 1341 -483 1375 389
rect -201 -542 1309 -508
<< locali >>
rect -270 424 -201 458
rect 1309 424 1375 458
rect -270 389 -236 424
rect -270 -508 -236 -483
rect 1341 389 1375 424
rect 1341 -508 1375 -483
rect -270 -542 -201 -508
rect 1309 -542 1375 -508
<< metal1 >>
rect -139 305 -80 392
rect 88 343 98 395
rect 190 343 200 395
rect 415 346 689 392
rect 904 343 914 395
rect 1006 343 1016 395
rect 1184 305 1242 392
rect -176 293 88 305
rect -176 117 -91 293
rect -39 117 88 293
rect -176 105 88 117
rect 200 105 360 305
rect 472 293 632 305
rect 459 117 469 293
rect 521 117 583 293
rect 635 117 645 293
rect 472 105 632 117
rect 744 105 904 305
rect 1016 293 1280 305
rect 1016 117 1143 293
rect 1195 117 1280 293
rect 1016 105 1280 117
rect 237 -18 324 105
rect 360 15 370 67
rect 462 15 472 67
rect 632 15 642 67
rect 734 15 744 67
rect 781 -18 869 105
rect 237 -69 869 -18
rect 89 -151 99 -99
rect 191 -151 201 -99
rect 237 -189 324 -69
rect 781 -189 869 -69
rect 905 -151 915 -99
rect 1007 -151 1017 -99
rect -174 -201 90 -189
rect -187 -377 -177 -201
rect -125 -377 90 -201
rect -174 -389 90 -377
rect 201 -389 361 -189
rect 473 -201 633 -189
rect 460 -377 470 -201
rect 522 -377 584 -201
rect 636 -377 646 -201
rect 473 -389 633 -377
rect 745 -389 905 -189
rect 1017 -201 1281 -189
rect 1017 -377 1232 -201
rect 1284 -377 1294 -201
rect 1017 -389 1281 -377
rect -136 -439 -78 -389
rect 361 -479 371 -427
rect 463 -430 473 -427
rect 633 -430 643 -427
rect 463 -475 643 -430
rect 463 -479 473 -475
rect 633 -479 643 -475
rect 735 -479 745 -427
rect 1185 -438 1243 -389
<< via1 >>
rect 98 343 190 395
rect 914 343 1006 395
rect -91 117 -39 293
rect 469 117 521 293
rect 583 117 635 293
rect 1143 117 1195 293
rect 370 15 462 67
rect 642 15 734 67
rect 99 -151 191 -99
rect 915 -151 1007 -99
rect -177 -377 -125 -201
rect 470 -377 522 -201
rect 584 -377 636 -201
rect 1232 -377 1284 -201
rect 371 -479 463 -427
rect 643 -479 735 -427
<< metal2 >>
rect 98 397 190 407
rect 0 367 31 368
rect -177 335 31 367
rect -177 -191 -130 335
rect -91 293 -39 303
rect -177 -201 -125 -191
rect -177 -387 -125 -377
rect -91 -430 -39 117
rect 0 64 31 335
rect 914 397 1006 407
rect 98 331 190 341
rect 251 346 521 392
rect 251 64 311 346
rect 469 293 521 346
rect 469 107 521 117
rect 583 346 856 392
rect 583 293 635 346
rect 583 107 635 117
rect 0 18 311 64
rect 370 67 462 77
rect 370 -18 462 15
rect 99 -69 462 -18
rect 642 67 734 77
rect 796 64 856 346
rect 914 331 1006 341
rect 1075 349 1284 385
rect 1075 64 1110 349
rect 796 18 1110 64
rect 1143 293 1195 303
rect 642 -18 734 15
rect 642 -69 1007 -18
rect 99 -99 191 -69
rect 915 -99 1007 -69
rect 99 -161 191 -151
rect 251 -148 522 -102
rect 251 -430 311 -148
rect 470 -201 522 -148
rect 470 -387 522 -377
rect 584 -148 856 -102
rect 584 -201 636 -148
rect 584 -387 636 -377
rect -91 -476 311 -430
rect 371 -425 463 -415
rect 371 -491 463 -481
rect 643 -425 735 -415
rect 796 -430 856 -148
rect 915 -161 1007 -151
rect 1143 -430 1195 117
rect 1232 -201 1284 349
rect 1232 -387 1284 -377
rect 796 -476 1195 -430
rect 643 -491 735 -481
<< via2 >>
rect 98 395 190 397
rect 98 343 190 395
rect 914 395 1006 397
rect 98 341 190 343
rect 914 343 1006 395
rect 914 341 1006 343
rect 371 -427 463 -425
rect 371 -479 463 -427
rect 371 -481 463 -479
rect 643 -427 735 -425
rect 643 -479 735 -427
rect 643 -481 735 -479
<< metal3 >>
rect 88 397 311 402
rect 88 341 98 397
rect 190 341 311 397
rect 88 336 311 341
rect 251 -420 311 336
rect 796 397 1016 402
rect 796 341 914 397
rect 1006 341 1016 397
rect 796 336 1016 341
rect 796 -420 856 336
rect 251 -425 473 -420
rect 251 -481 371 -425
rect 463 -481 473 -425
rect 251 -486 473 -481
rect 633 -425 856 -420
rect 633 -481 643 -425
rect 735 -481 856 -425
rect 633 -486 856 -481
use sky130_fd_pr__pfet_01v8_BH5GQ5  sky130_fd_pr__pfet_01v8_BH5GQ5_0
timestamp 1729185150
transform 1 0 552 0 1 205
box -552 -200 552 200
use sky130_fd_pr__pfet_01v8_BH5GQ5  sky130_fd_pr__pfet_01v8_BH5GQ5_1
timestamp 1729185150
transform 1 0 553 0 1 -289
box -552 -200 552 200
use sky130_fd_pr__pfet_01v8_LA8JHL  sky130_fd_pr__pfet_01v8_LA8JHL_0
timestamp 1729187732
transform 1 0 -109 0 1 -325
box -109 -164 109 198
use sky130_fd_pr__pfet_01v8_LA8JHL  sky130_fd_pr__pfet_01v8_LA8JHL_1
timestamp 1729187732
transform 1 0 1214 0 1 -325
box -109 -164 109 198
use sky130_fd_pr__pfet_01v8_MA8JHN  sky130_fd_pr__pfet_01v8_MA8JHN_0
timestamp 1729187732
transform 1 0 -109 0 1 241
box -109 -198 109 164
use sky130_fd_pr__pfet_01v8_MA8JHN  sky130_fd_pr__pfet_01v8_MA8JHN_1
timestamp 1729187732
transform 1 0 1213 0 1 241
box -109 -198 109 164
<< labels >>
flabel metal3 224 367 224 367 0 FreeSans 160 0 0 0 VIN
port 0 nsew
flabel metal2 216 -46 216 -46 0 FreeSans 160 0 0 0 VIP
port 1 nsew
flabel metal1 552 -44 552 -44 0 FreeSans 160 0 0 0 D5
port 2 nsew
flabel metal2 1258 -47 1259 -46 0 FreeSans 160 0 0 0 OUT
port 3 nsew
flabel nsubdiffcont 553 439 553 439 0 FreeSans 160 0 0 0 VDD
port 4 nsew
flabel metal2 1171 -51 1171 -51 0 FreeSans 160 0 0 0 D6
port 5 nsew
<< end >>
