magic
tech sky130A
magscale 1 2
timestamp 1729187732
<< error_p >>
rect -29 145 29 151
rect -29 111 -17 145
rect -29 105 29 111
<< nwell >>
rect -109 -198 109 164
<< pmos >>
rect -15 -136 15 64
<< pdiff >>
rect -73 52 -15 64
rect -73 -124 -61 52
rect -27 -124 -15 52
rect -73 -136 -15 -124
rect 15 52 73 64
rect 15 -124 27 52
rect 61 -124 73 52
rect 15 -136 73 -124
<< pdiffc >>
rect -61 -124 -27 52
rect 27 -124 61 52
<< poly >>
rect -33 145 33 161
rect -33 111 -17 145
rect 17 111 33 145
rect -33 95 33 111
rect -15 64 15 95
rect -15 -162 15 -136
<< polycont >>
rect -17 111 17 145
<< locali >>
rect -33 111 -17 145
rect 17 111 33 145
rect -61 52 -27 68
rect -61 -140 -27 -124
rect 27 52 61 68
rect 27 -140 61 -124
<< viali >>
rect -17 111 17 145
rect -61 -124 -27 52
rect 27 -124 61 52
<< metal1 >>
rect -29 145 29 151
rect -29 111 -17 145
rect 17 111 29 145
rect -29 105 29 111
rect -67 52 -21 64
rect -67 -124 -61 52
rect -27 -124 -21 52
rect -67 -136 -21 -124
rect 21 52 67 64
rect 21 -124 27 52
rect 61 -124 67 52
rect 21 -136 67 -124
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
