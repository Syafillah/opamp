magic
tech sky130A
magscale 1 2
timestamp 1729362362
<< viali >>
rect 1353 2802 1387 2836
rect 2378 717 2414 751
<< metal1 >>
rect 2152 3094 2198 3140
rect 811 2836 1399 2842
rect 811 2802 1353 2836
rect 1387 2802 1399 2836
rect 811 2797 1399 2802
rect 1341 2796 1399 2797
rect 1113 2678 1945 2733
rect 1115 1561 1183 2678
rect 1654 2367 1664 2547
rect 1716 2367 1726 2547
rect 2451 1851 2461 1903
rect 2548 1851 2558 1903
rect 1105 1509 1115 1561
rect 1183 1509 1193 1561
rect 828 905 862 947
rect 1910 905 2078 906
rect 819 835 2078 905
rect 828 834 862 835
rect 1910 629 2078 835
rect 2366 751 2426 1032
rect 2366 717 2378 751
rect 2414 717 2426 751
rect 2366 710 2426 717
rect 2683 619 2740 675
rect 547 111 557 163
rect 699 111 709 163
<< via1 >>
rect 1664 2367 1716 2547
rect 2461 1851 2548 1903
rect 1115 1509 1183 1561
rect 557 111 699 163
<< metal2 >>
rect 1662 2547 1718 2557
rect 1662 2357 1718 2367
rect 2686 2144 2762 2318
rect 2460 2084 2762 2144
rect 2460 2075 2761 2084
rect 2461 1903 2548 2075
rect 2461 1841 2548 1851
rect 820 1561 1183 1571
rect 820 1509 1115 1561
rect 820 1500 1183 1509
rect 1115 1499 1183 1500
rect 1153 845 2256 892
rect 557 163 699 173
rect 1153 163 1259 845
rect 2211 570 2256 845
rect 547 111 557 163
rect 699 111 1259 163
rect 547 103 1259 111
rect 547 102 1162 103
rect 557 101 699 102
<< via2 >>
rect 1662 2367 1664 2547
rect 1664 2367 1716 2547
rect 1716 2367 1718 2547
<< metal3 >>
rect 1711 3084 1823 3155
rect 1652 2547 1728 2552
rect 1652 2367 1662 2547
rect 1718 2367 1728 2547
rect 1652 2362 1728 2367
rect 1660 2129 1720 2362
rect 1660 2043 2207 2129
rect 2147 1785 2207 2043
use nmos_diffamp  nmos_diffamp_0
timestamp 1729221670
transform 1 0 1712 0 1 1498
box -324 -536 1254 512
use nmoscs  nmoscs_0
timestamp 1729233261
transform 1 0 1836 0 1 109
box -384 -798 1072 677
use pmocs  pmocs_0
timestamp 1729233261
transform 1 0 184 0 1 877
box -184 -877 814 1995
use pmos_diffamp  pmos_diffamp_0
timestamp 1729213131
transform 1 0 1623 0 1 2748
box -306 -578 1411 494
<< labels >>
flabel metal1 1158 2820 1158 2820 0 FreeSans 800 0 0 0 VDD
port 0 nsew
flabel metal3 1929 2091 1929 2091 0 FreeSans 800 0 0 0 OUT
port 1 nsew
flabel metal1 2397 912 2397 912 0 FreeSans 800 0 0 0 GND
port 2 nsew
flabel metal1 2711 652 2711 652 0 FreeSans 800 0 0 0 RS
port 3 nsew
flabel metal1 2176 3120 2176 3120 0 FreeSans 800 0 0 0 VIP
port 4 nsew
flabel metal3 1769 3120 1769 3120 0 FreeSans 800 0 0 0 VIN
port 5 nsew
<< end >>
